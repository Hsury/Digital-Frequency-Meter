LIBRARY IEEE; --数字频率计
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY FREQTEST IS
	PORT (CLK : IN STD_LOGIC; --50MHz标准频率时钟
         FSIN : IN STD_LOGIC; --待测频率
         DUAN : OUT STD_LOGIC_VECTOR (7 DOWNTO 0); --数码管段
			WEI : OUT STD_LOGIC_VECTOR (5 DOWNTO 0)); --数码管位
END FREQTEST;
ARCHITECTURE struc OF FREQTEST IS
	COMPONENT DIVFREQ
	PORT(FSTD : IN STD_LOGIC;
	     CLKBUS : OUT STD_LOGIC_VECTOR (8 DOWNTO 0));
	END COMPONENT;
	COMPONENT TESTCTL
	PORT(CLK : IN STD_LOGIC;
	     TSTEN : OUT STD_LOGIC;
		  CLR_CNT : OUT STD_LOGIC;
		  Load : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT CNT10
	PORT(CLK : IN STD_LOGIC;
	     CLR : IN STD_LOGIC;
		  ENA : IN STD_LOGIC;
		  CQ : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		  CARRY_OUT : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT REG24B
	PORT (Load : IN STD_LOGIC;
	      DIN : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			DOUT : OUT STD_LOGIC_VECTOR (23 DOWNTO 0));
	END COMPONENT;
	COMPONENT LEDCTRL
	PORT(CLK : IN STD_LOGIC;
	     DATA : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
	     CURSOR : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		  NUM : OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
	END COMPONENT;
	COMPONENT DECODER3TO8
	PORT(BIN3BIT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	     WEI : OUT STD_LOGIC_VECTOR (5 DOWNTO 0));
	END COMPONENT;
	COMPONENT SEG8
	PORT(DATA : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     DOT : IN STD_LOGIC;
	     DUAN : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
	END COMPONENT;
	SIGNAL CLKBUS : STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL Load1, TSTEN1, CLR_CNT1 : STD_LOGIC;
	SIGNAL DTO1 : STD_LOGIC_VECTOR (23 DOWNTO 0);
	SIGNAL CARRY_OUT1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL DOUT : STD_LOGIC_VECTOR (23 DOWNTO 0);
	SIGNAL BIN3BIT : STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL NUM : STD_LOGIC_VECTOR (3 DOWNTO 0);
BEGIN
	U0 : DIVFREQ PORT MAP(FSTD => CLK,
	                      CLKBUS => CLKBUS);
	U1 : TESTCTL PORT MAP(CLK => CLKBUS(1),
	                      TSTEN => TSTEN1,
								 CLR_CNT => CLR_CNT1,
								 Load => Load1);
	U2 : REG24B PORT MAP(Load => Load1,
	                     DIN => DTO1,
								DOUT => DOUT);
	U3 : CNT10 PORT MAP(CLK => CLKBUS(6), --待测频率在这里传入
	                    CLR => CLR_CNT1,
							  ENA => TSTEN1,
							  CQ => DTO1(3 DOWNTO 0),
							  CARRY_OUT => CARRY_OUT1(0));
	U4 : CNT10 PORT MAP(CLK => CARRY_OUT1(0),
	                    CLR => CLR_CNT1,
							  ENA => TSTEN1,
							  CQ => DTO1(7 DOWNTO 4),
							  CARRY_OUT => CARRY_OUT1(1));
	U5 : CNT10 PORT MAP(CLK => CARRY_OUT1(1),
	                    CLR => CLR_CNT1,
							  ENA => TSTEN1,
							  CQ => DTO1(11 DOWNTO 8),
	                    CARRY_OUT => CARRY_OUT1(2));
	U6 : CNT10 PORT MAP(CLK => CARRY_OUT1(2),
	                    CLR => CLR_CNT1,
	                    ENA => TSTEN1,
							  CQ => DTO1(15 DOWNTO 12),
	                    CARRY_OUT => CARRY_OUT1(3));
	U7 : CNT10 PORT MAP(CLK => CARRY_OUT1(3),
	                    CLR => CLR_CNT1,
							  ENA => TSTEN1,
							  CQ => DTO1(19 DOWNTO 16),
	                    CARRY_OUT => CARRY_OUT1(4));
	U8 : CNT10 PORT MAP(CLK => CARRY_OUT1(4),
	                    CLR => CLR_CNT1,
							  ENA => TSTEN1,
							  CQ => DTO1(23 DOWNTO 20));
	U9 : LEDCTRL PORT MAP(CLK => CLKBUS(4), --设置数码管刷新频率为1KHz
	                      DATA => DOUT,
								 CURSOR => BIN3BIT,
								 NUM => NUM);
	U10 : DECODER3TO8 PORT MAP(BIN3BIT => BIN3BIT,
	                           WEI => WEI);
	U11 : SEG8 PORT MAP(DATA => NUM,
	                    DOT => '0',
							  DUAN => DUAN);
END struc;