LIBRARY IEEE; --测频控制信号发生器
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY TESTCTL IS
	PORT (CLK : IN STD_LOGIC; --1Hz测频控制时钟
         TSTEN : OUT STD_LOGIC; --计数器时钟使能
         CLR_CNT : OUT STD_LOGIC; --计数器清零
         Load : OUT STD_LOGIC); --输出锁存信号
END TESTCTL;
ARCHITECTURE behav OF TESTCTL IS
	SIGNAL Div2CLK : STD_LOGIC;
BEGIN
	PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK='1' THEN --1Hz时钟二分频
			Div2CLK<=NOT Div2CLK;
		END IF;
	END PROCESS;
	PROCESS(CLK, Div2CLK)
	BEGIN
		IF CLK='0' AND Div2CLK='0' THEN
			CLR_CNT<='1'; --产生计数器清零信号
		ELSE
			CLR_CNT<='0';
		END IF;
	END PROCESS;
	Load<=NOT Div2CLK;
	TSTEN<=CLK;
END behav;