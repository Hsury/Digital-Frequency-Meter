LIBRARY IEEE; --10进制9级分频器
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DIVFREQ IS
	PORT(FSTD : IN STD_LOGIC;
	     CLKBUS : OUT STD_LOGIC_VECTOR (8 DOWNTO 0)); --映射10MHz到0.1Hz
END DIVFREQ;
ARCHITECTURE behav OF DIVFREQ IS
	SIGNAL CO0, CO1, CO2, CO3, CO4, CO5, CO6, CO7, CO8 : STD_LOGIC;
BEGIN
	PROCESS (FSTD)
		VARIABLE CNT0 : INTEGER RANGE 0 TO 4;
	BEGIN
		IF RISING_EDGE(FSTD) THEN
			IF CNT0<2 THEN
				CO0<='1';
				CNT0:=CNT0+1;
			ELSIF CNT0<4 THEN
				CO0<='0';
				CNT0:=CNT0+1;
			ELSE
				CNT0:=0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (CO0)
		VARIABLE CNT1 : INTEGER RANGE 0 TO 9;
	BEGIN
		IF RISING_EDGE(CO0) THEN
			IF CNT1<5 THEN
				CO1<='1';
				CNT1:=CNT1+1;
			ELSIF CNT1<9 THEN
				CO1<='0';
				CNT1:=CNT1+1;
			ELSE
				CNT1:=0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (CO1)
		VARIABLE CNT2 : INTEGER RANGE 0 TO 9;
	BEGIN
		IF RISING_EDGE(CO1) THEN
			IF CNT2<5 THEN
				CO2<='1';
				CNT2:=CNT2+1;
			ELSIF CNT2<9 THEN
				CO2<='0';
				CNT2:=CNT2+1;
			ELSE
				CNT2:=0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (CO2)
		VARIABLE CNT3 : INTEGER RANGE 0 TO 9;
	BEGIN
		IF RISING_EDGE(CO2) THEN
			IF CNT3<5 THEN
				CO3<='1';
				CNT3:=CNT3+1;
			ELSIF CNT3<9 THEN
				CO3<='0';
				CNT3:=CNT3+1;
			ELSE
				CNT3:=0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (CO3)
		VARIABLE CNT4 : INTEGER RANGE 0 TO 9;
	BEGIN
		IF RISING_EDGE(CO3) THEN
			IF CNT4<5 THEN
				CO4<='1';
				CNT4:=CNT4+1;
			ELSIF CNT4<9 THEN
				CO4<='0';
				CNT4:=CNT4+1;
			ELSE
				CNT4:=0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (CO4)
		VARIABLE CNT5 : INTEGER RANGE 0 TO 9;
	BEGIN
		IF RISING_EDGE(CO4) THEN
			IF CNT5<5 THEN
				CO5<='1';
				CNT5:=CNT5+1;
			ELSIF CNT5<9 THEN
				CO5<='0';
				CNT5:=CNT5+1;
			ELSE
				CNT5:=0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (CO5)
		VARIABLE CNT6 : INTEGER RANGE 0 TO 9;
	BEGIN
		IF RISING_EDGE(CO5) THEN
			IF CNT6<5 THEN
				CO6<='1';
				CNT6:=CNT6+1;
			ELSIF CNT6<9 THEN
				CO6<='0';
				CNT6:=CNT6+1;
			ELSE
				CNT6:=0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (CO6)
		VARIABLE CNT7 : INTEGER RANGE 0 TO 9;
	BEGIN
		IF RISING_EDGE(CO6) THEN
			IF CNT7<5 THEN
				CO7<='1';
				CNT7:=CNT7+1;
			ELSIF CNT7<9 THEN
				CO7<='0';
				CNT7:=CNT7+1;
			ELSE
				CNT7:=0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (CO7)
		VARIABLE CNT8 : INTEGER RANGE 0 TO 9;
	BEGIN
		IF RISING_EDGE(CO7) THEN
			IF CNT8<5 THEN
				CO8<='1';
				CNT8:=CNT8+1;
			ELSIF CNT8<9 THEN
				CO8<='0';
				CNT8:=CNT8+1;
			ELSE
				CNT8:=0;
			END IF;
		END IF;
	END PROCESS;
	CLKBUS<=CO0 & CO1 & CO2 & CO3 & CO4 & CO5 & CO6 & CO7 & CO8;
END behav;