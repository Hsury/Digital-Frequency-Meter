LIBRARY IEEE; --3-8译码器(数码管位选控制器)
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DECODER3TO8 IS
	PORT(BIN3BIT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	     WEI : OUT BIT_VECTOR (5 DOWNTO 0));
END DECODER3TO8;
ARCHITECTURE behav OF DECODER3TO8 IS
BEGIN
	WEI<="011111" ROR CONV_INTEGER(BIN3BIT);
END behav;