LIBRARY IEEE; --24 位锁存器
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY REG24B IS
	PORT (Load : IN STD_LOGIC;
         DIN : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
         DOUT : OUT STD_LOGIC_VECTOR (23 DOWNTO 0));
END REG24B;
ARCHITECTURE behav OF REG24B IS
BEGIN
		PROCESS(Load, DIN)
		BEGIN
			IF Load'EVENT AND Load='1' THEN
				DOUT<=DIN; --锁存输入数据
			END IF;
		END PROCESS;
END behav;