--主控制器模块 2017/05/23
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CTRL IS
	PORT (CLK_SYNC : IN STD_LOGIC;	--同步信号
	      CREG : BUFFER STD_LOGIC;	--锁存信号
	      CLR : OUT STD_LOGIC;	--清零信号
	      CP : OUT STD_LOGIC);	--计数使能信号
END CTRL;

ARCHITECTURE BEHAV OF CTRL IS
	SIGNAL C : STD_LOGIC;
BEGIN
	PROCESS (CLK_SYNC)
	BEGIN
		IF RISING_EDGE(CLK_SYNC) THEN
			C <= NOT C;
		END IF;
	END PROCESS;
	
	PROCESS (C, CLK_SYNC)
	BEGIN
		IF C = '0' AND CLK_SYNC = '0' THEN
			CLR <= '1';
		ELSE
			CLR <= '0';
		END IF;
	END PROCESS;
	
	CREG <= NOT C;
	CP <= C;
END BEHAV;